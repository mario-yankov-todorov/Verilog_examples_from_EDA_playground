/*
*	M. Todorov 2021
*/

`timescale 1ns / 1ps

module code_lock
 	(
		input 	A,
		input 	M,
		input 	C,
		
		output	F
  	);
  
  	assign F = M | (A & C);
  
endmodule
