interface intf(input logic clk, rst);
	
		// Declare the signals
		logic 			button;
		logic  [8	-1:0] 	valid_in;
	
endinterface